-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Tue Nov 22 00:09:01 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PARTE_D IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        Z3 : OUT STD_LOGIC;
        Z2 : OUT STD_LOGIC;
        Z1 : OUT STD_LOGIC;
        Z0 : OUT STD_LOGIC
    );
END PARTE_D;

ARCHITECTURE BEHAVIOR OF PARTE_D IS
    TYPE type_fstate IS (E,F,G,C,D,A,B);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= B;
            Z3 <= '0';
            Z2 <= '0';
            Z1 <= '0';
            Z0 <= '0';
        ELSE
            Z3 <= '0';
            Z2 <= '0';
            Z1 <= '0';
            Z0 <= '0';
            CASE fstate IS
                WHEN E =>
                    reg_fstate <= F;

                    Z0 <= '0';

                    Z1 <= '1';

                    Z3 <= '0';

                    Z2 <= '1';
                WHEN F =>
                    IF ((x = '0')) THEN
                        reg_fstate <= G;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= D;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= F;
                    END IF;

                    Z0 <= '1';

                    Z1 <= '1';

                    Z3 <= '1';

                    Z2 <= '1';
                WHEN G =>
                    reg_fstate <= A;

                    Z0 <= '1';

                    Z1 <= '0';

                    Z3 <= '1';

                    Z2 <= '0';
                WHEN C =>
                    reg_fstate <= D;

                    Z0 <= '0';

                    Z1 <= '0';

                    Z3 <= '1';

                    Z2 <= '1';
                WHEN D =>
                    reg_fstate <= A;

                    Z0 <= '0';

                    Z1 <= '1';

                    Z3 <= '1';

                    Z2 <= '1';
                WHEN A =>
                    IF ((x = '0')) THEN
                        reg_fstate <= E;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    Z0 <= '0';

                    Z1 <= '0';

                    Z3 <= '0';

                    Z2 <= '0';
                WHEN B =>
                    reg_fstate <= C;

                    Z0 <= '0';

                    Z1 <= '0';

                    Z3 <= '1';

                    Z2 <= '0';
                WHEN OTHERS => 
                    Z3 <= 'X';
                    Z2 <= 'X';
                    Z1 <= 'X';
                    Z0 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
